--LED灯控制模块--
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY LED IS
   PORT(GC_MODE,SW_MODE:IN INTEGER RANGE 0 TO 2;         --过程选择和水位选择信号--
	     SET:IN INTEGER RANGE 0 TO 3;               		--模式选择信号--
	     GC_L,SW_L:OUT STD_LOGIC_VECTOR(2 DOWNTO 0);      --过程和水位输出LED灯信号（3个灯）--
		  MS_L:OUT STD_LOGIC_VECTOR(3 DOWNTO 0));          --模式输出LED灯信号（4个灯）--
END ENTITY LED;

ARCHITECTURE L OF LED IS
BEGIN 
p:PROCESS(GC_MODE,SW_MODE,SET)
BEGIN
--过程指示灯部分--
IF(GC_MODE=0)THEN  GC_L<="100";
ELSIF(GC_MODE=1)THEN  GC_L<="010";
ELSIF(GC_MODE=2)THEN  GC_L<="001";
ELSE NULL;
END IF;
--水位指示灯部分--
IF(SW_MODE=0)THEN  SW_L<="100";
ELSIF(SW_MODE=1)THEN  SW_L<="010";
ELSIF(SW_MODE=2)THEN  SW_L<="001";
ELSE NULL;
END IF;
--模式指示灯部分--
IF(SET=0)THEN  MS_L<="1000";
ELSIF(SET=1)THEN  MS_L<="0100";
ELSIF(SET=2)THEN  MS_L<="0010";
ELSIF(SET=3)THEN  MS_L<="0001";
ELSE NULL;
END IF;
END PROCESS p;
END ARCHITECTURE L;